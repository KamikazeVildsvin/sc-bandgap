** sch_path:
*+ /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/sc-bandgap/test-tg.sch
**.subckt test-tg
V1 VDD VSS 1.8
V2 VSS 0 0
x1 GATEP DRAIN SOURCE GATEN VDD VSS transmissiongate WP=1u LP=0.26u WN=0.26u LN=0.26u m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  transmissiongate.sym # of pins=4
** sym_path:
*+ /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/sc-bandgap/transmissiongate.sym
** sch_path:
*+ /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/sc-bandgap/transmissiongate.sch
.subckt transmissiongate  GP DPIN SPIN GN  VDDBPIN  VSSBPIN   WP=1u LP=0.26u WN=0.26u LN=0.26u
*.iopin DPIN
*.iopin SPIN
*.iopin GN
*.iopin GP
XM1 DPIN GN SPIN VSSBPIN sky130_fd_pr__nfet_01v8 L=LN W=WN nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=M m=M
XM2 DPIN GP SPIN VDDBPIN sky130_fd_pr__pfet_01v8 L=LP W=WP nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=M m=M
.ends

.end
