** sch_path:
*+ /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/sc-bandgap/sc_bandgap.sch
**.subckt sc_bandgap VDD VREF VSS
*.iopin VDD
*.opin VREF
*.iopin VSS
I2 VDD VBE2 10u
I1 VDD VBE1 10u
XQ1 VSS VSS VBE1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=10
XQ2 VSS VSS VBE2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
V1 VDD VSS 1.8
.save i(v1)
V2 CLK VSS PULSE(0 1.8 0 {t_rise} {t_fall} {(1-dutycycle)*1/clk_freq} {1/clk_freq} 0)
.save i(v2)
V4 VSS 0 0
.save i(v4)
XC1K CAP1K X sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=4*9 m=4*9
XC1 CAP1 X sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=4 m=4
XC3 CAP3 VREF sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=6 m=6
XC2 X CAP2 sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=4*2 m=4*2
XM1 CAP1 PHI2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.26 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 CAP3 PHI1 X VSS sky130_fd_pr__nfet_01v8 L=0.26 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 CAP3 PHI2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.26 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 CAP2 PHI1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.26 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
x1 N_PHI2 VBE1 CAP1K PHI2 VDD VSS transmissiongate W_P=2 L_P=0.26 W_N=1 L_N=0.26 m=1
x2 N_PHI1 VBE2 CAP1K PHI1 VDD VSS transmissiongate W_P=2 L_P=0.26 W_N=1 L_N=0.26 m=1
x3 N_PHI1 VBE2 CAP1 PHI1 VDD VSS transmissiongate W_P=2 L_P=0.26 W_N=1 L_N=0.26 m=1
.save v(vbe2)
.save v(vbe1)
x8 CLK net1 net3 VDD VSS lvnand WidthN=1 LenN=0.15 WidthP=1 LenP=0.15 m=1
x9 net4 net2 net5 VDD VSS lvnand WidthN=1 LenN=0.15 WidthP=1 LenP=0.15 m=1
x10 net4 CLK VDD VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x11 PHI2 net2 VDD VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x12 net6 net3 VDD VSS not W_N=0.5 L_N=1 W_P=1 L_P=1 m=1
x13 net7 net6 VDD VSS not W_N=0.5 L_N=1 W_P=1 L_P=1 m=1
x14 net8 net7 VDD VSS not W_N=0.5 L_N=1 W_P=1 L_P=1 m=1
x15 net2 net8 VDD VSS not W_N=0.5 L_N=1 W_P=1 L_P=1 m=1
x16 net9 net5 VDD VSS not W_N=0.5 L_N=1 W_P=1 L_P=1 m=1
x17 net10 net9 VDD VSS not W_N=0.5 L_N=1 W_P=1 L_P=1 m=1
x18 net11 net10 VDD VSS not W_N=0.5 L_N=1 W_P=1 L_P=1 m=1
x19 net1 net11 VDD VSS not W_N=0.5 L_N=1 W_P=1 L_P=1 m=1
x20 PHI1 net1 VDD VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x22 N_PHI1 PHI1 VDD VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x4 N_PHI2 PHI2 VDD VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x5 N_PHI2 CAP2 VREF PHI2 VDD VSS transmissiongate W_P=2 L_P=0.26 W_N=1 L_N=0.26 m=1
x6 VSS VREF X VDD VSS opamp_onepole gain=1e4 f3db=2e6
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



* Parameters *
.param clk_freq = 1Meg
.param dutycycle = 0.5
.param t_rise = 1n
.param t_fall = 1n

* Switch model *
.model SWITCH1 sw vt=1 vh=0.2 ron=1k roff=1Meg

* Options *
.options wnflag=1 RELTOL=0.001
*.options wnflag=1 METHOD=GEAR ITL4=100 CHGTOL=1e-15 TRTOL=1 RELTOL=0.0001 VNTOL=0.1u
.options savecurrents
.save all
.save @m.xm1.msky130_fd_pr__nfet_01v8[gds]
.save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
.save @m.xm2.msky130_fd_pr__nfet_01v8[gds]
.save @q.xq1.qsky130_fd_pr__pnp_05v5_W3p40L3p40[p]

* Control *
.control
let run = 1
set temp=0
while run <= 3
   if run > 1
      reset
      set appendwrite
   end
   let dtemp = 0 + 40*(run-1)
   set temp=$&dtemp
   tran 1n 10u 8u
   write sc_bandgap.raw
   let run = run + 1
end
reset
op
set appendwrite
write sc_bandgap.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  transmissiongate.sym # of pins=4
** sym_path:
*+ /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/sc-bandgap/transmissiongate.sym
** sch_path:
*+ /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/sc-bandgap/transmissiongate.sch
.subckt transmissiongate GP DPIN SPIN GN  VDDBPIN  VSSBPIN   W_P=1 L_P=0.2 W_N=1 L_N=0.2
*.iopin DPIN
*.iopin SPIN
*.ipin GP
*.ipin GN
XM1 DPIN GN SPIN VSSBPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=m m=m
XM2 DPIN GP SPIN VDDBPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=m m=m
.ends


* expanding   symbol:  sky130_tests/lvnand.sym # of pins=3
** sym_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/lvnand.sym
** sch_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/lvnand.sch
.subckt lvnand A B Y  VCCPIN  VSSPIN   WidthN=1 LenN=0.15 WidthP=1 LenP=0.15
*.ipin A
*.ipin B
*.opin Y
XM1 Y B S VSSPIN sky130_fd_pr__nfet_01v8 L=LenN W=WidthN nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=LenP W=WidthP nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y B VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=LenP W=WidthP nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 S A VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=LenN W=WidthN nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sky130_tests/not.sym # of pins=2
** sym_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sym
** sch_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sch
.subckt not y a  VCCPIN  VSSPIN      W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  opamp_onepole.sym # of pins=3
** sym_path:
*+ /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/sc-bandgap/opamp_onepole.sym
** sch_path:
*+ /Users/nlv/Documents/DTU/9.Semester/IC-Open-Source/xschem-projects/sc-bandgap/opamp_onepole.sch
.subckt opamp_onepole POS OUT NEG  VDDPIN  VSSPIN   gain=1e4 f3db=2e6
*.opin OUT
*.ipin POS
*.ipin NEG
E1 VDIFF VSSPIN VOL=' (V(POS)-V(NEG))*gain > V(VDDPIN) ? V(VDDPIN) : (V(POS)-V(NEG))*gain < V(VSSPIN) ? V(VSSPIN) : (V(POS)-V(NEG))*gain '
R3 SR VDIFF 1k m=1
C2 SR VSSPIN {1/(2*3.149*1e3*f3db)} m=1
E2 OUT VSSPIN VOL=' V(SR)*1 '
.ends

.end
